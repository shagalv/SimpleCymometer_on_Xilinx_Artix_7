
module oled_clear(
    input send_done,
    output reg spi_send,
    output reg[7:0] spi_data,
    input clk,
    output dc,
    input clear_start,
    output clear_done,
    input reset

);
    reg [3:0]cur_st,nxt_st;
    assign dc=(cur_st==4)?1:0;
    assign clear_done=(cur_st==6)?1:0;
    //assign spi_send=(cur_st==1 | 2 | 3 | 4)?1:0;

    reg [7:0]x_tmp,y_tmp;  
    wire [7:0]     Set_pos_0=8'hb0 | y_tmp,
                    Set_pos_1= (x_tmp[7:4] & 4'hf) | 8'h10,
                    Set_pos_2= (x_tmp[3:0] & 4'hf);
    
    reg [47:0]write_data_tmp;
    reg [3:0]count;
    
    
    always@(posedge clk or posedge reset)
        if(reset)
            cur_st<=0;
        else if(cur_st==1 | cur_st==2 | cur_st==3 | cur_st==4 ) 
           begin if(send_done)  cur_st<=nxt_st; end
        else cur_st<=nxt_st;

    always@(*)
    begin
        nxt_st=cur_st;
        case(cur_st)
            0:begin if(clear_start)                 nxt_st=cur_st+1; end
            1:begin            nxt_st=cur_st+1; end
            2:begin            nxt_st=cur_st+1; end
            3:begin            nxt_st=cur_st+1; end
            4:begin            nxt_st=cur_st+1; end  
            5:if(x_tmp==127 && y_tmp==7) begin nxt_st=6;         end
              else  begin               nxt_st=1;        end  
            6:begin                     nxt_st=0;        end
            default:begin nxt_st=0;end
        endcase
    end
    
    always@(*)
        if(reset)
        begin
            spi_data=0;
            spi_send=0;
        end
        else case(cur_st)
            0:begin spi_data = 0;                      spi_send=0;    end 
            1:begin spi_data = Set_pos_0;              spi_send=1;    end
            2:begin spi_data = Set_pos_1;              spi_send=1;    end
            3:begin spi_data = Set_pos_2;              spi_send=1;    end      
            4:begin spi_data = 0;                      spi_send=1;    end
            5:spi_send=0;
            endcase
       
    always@(posedge clk or posedge reset)
        if(reset)
        begin
            x_tmp<=0;
            y_tmp<=0;
            write_data_tmp<=0;
            count<=0;
        end
        else case(cur_st)
            0:begin
                x_tmp<=0;
                y_tmp<=0;
                count<=0;
              end
            5:begin
                //if(x_tmp>122) y_tmp<=y_tmp+1;
                if(x_tmp==130)
                begin
                     y_tmp<=y_tmp+1;
                     x_tmp<=0;
                end
                else x_tmp<=x_tmp+1;
              end
        endcase

 endmodule
